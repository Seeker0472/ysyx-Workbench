module example(
  input a,
  input b,
  // input clk,
  output f
);
  assign f = a ^ b;
endmodule
